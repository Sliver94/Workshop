* ADG1421 SPICE Macro-model
* Generic Desc: 2.1 O On Resistance, �15 V/+12 V/�5 V iCMOS Dual SPST Switches
* Developed by: MPorley / ADGT
* Revision History: 1.0 (11/2019)
* Copyright 2019 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* Begin Notes:
* The model will work on Vdd/Vss from 5V to 16.5V single supply and +/-4.5V to +/-16.5V dual supply.
* The model provides parametric specifications at +/-16.5V only and is not variable with Vdd and Vss changes. Please see datasheet page 3. 
* The model is operational at RESET/VL level from V and 15V only. 
* Ensure 120us from the time of power-up or RESET before any logic command is issued. 
*
* Not Modeled:
* SPI Line interface and functionality is not modeled.
* The model would instead use a parallel line interface to control the switches.
* Please see Connections Section below.
*
* Parameters modeled include:
*	On Resistance
*	Ton and Toff
*	Break-Before-Make
*	Off Isolation
*	Crosstalk
*	Supply Currents: Iss/Idd
*	Bandwidth
*	Charge Injection
* Connections
*      1  = S1
*      2  = S2
*      3  = NC
*      4  = GND
*      5  = VDD
*      6  = IN2
*      7  = IN1
*      8  = VSS
*      9  = D2
*      10  = D1
*
.SUBCKT ADG1421 1 2 4 5 6 7 8 9 10

.MODEL VON VSWITCH(Von=5 Voff=0.8 Ron=0.001 Roff=1000000000000)
.MODEL VEN VSWITCH(Von=5 Voff=0.8 Ron=135000 Roff=215000)
.MODEL VRESET VSWITCH(Von=5 Voff=0.8 Ron= Roff=)
.MODEL DCLAMP D(IS=1E-15 IBV=1E-13)


* CROSSTALK
C12X 1 2 0.6E-012

* IDD/ISS
I1 5 4 0.002E-006
I2 8 4 0.002E-006

* Configuration: SPST 2:2 
 
 
** SWITCH 1 **
*
* ESD PROTECTION DIODES
D11 8 10 DCLAMP
D12 10 5 DCLAMP
D13 8 1 DCLAMP
D14 1 5 DCLAMP
*
* OFF ISOLATION
C11 1 10 1.9E-012
*
* CHARGE INJECTION
C12 10 140 2E-012
C13 1 140 2E-012
*
* CD/CS OFF AND BANDWIDTH
C14 1 4 12E-012
C15 10 4 15e-012
*
* ON RESISTANCE
Ech155 1555 4 VALUE = { IF ((ABS(V(1)))>(ABS(V(184))),V(1),V(10)) }
R155 1555 4 1G
R11 137 10 0.001
S111 136 141 1141 4 VON
Ech111 1141 4 VALUE = { IF (V(1555)<-13.5,5,0) }
Ech11 141 4 VALUE = { IF (V(1555)<-13.5,1.66666666666668E-02*(V(1555)--13.5)+2.45,0) }
S112 136 146 1146 4 VON
Ech112 1146 4 VALUE = { IF ((V(1555)>=-13.5) & (V(1555)<=13.5),5,0) }
Ech12 146 4 VALUE = { IF ((V(1555)>=-13.5) & (V(1555)<=13.5),((2.45-1.7)/((-13.5--0.796884641094606)*(-13.5--0.796884641094606)))*(V(1555)--0.796884641094606)*(V(1555)--0.796884641094606) + 1.7,0) }
S113 136 144 1144 4 VON
Ech113 1144 4 VALUE = { IF (V(1555)>13.5,5,0) }
Ech13 144 4 VALUE = { IF (V(1555)>13.5,-1.66666666666666E-02*(V(1555)-13.5)+2.65,0) }
RIN1	136 4	1G
EOUT1 137 181	POLY(2) (136,4) (180,4) 0 0 0 0 0.999/1000
FCOPY1	4 180 VSENSE1 1
RSENSOR1 180 4	1K
VSENSE1 181 184	0
*
* TON/ TOFF/ BBM
S11 182 184 140 4 VON
S12 143 138 143 4 VEN
Ech14 143 4 VALUE = { IF(V(7)>=2.0, 5 , 0.8 ) }
eV1 140 4 138 4 1
C16 138 4 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S13 1 182 185 4 VON
S14 142 185 142 4 VON
Ech15 142 4 VALUE = { IF((V(8)<=-0.5 & V(8)>=-16.5) & (V(5)<=16.5 & V(5)>=4.5), 5 , 0.01 ) }
S15 139 185 139 4 VON
Ech16 139 4 VALUE = { IF((V(8)>=-0.5 & (V(5)<=16.5 & V(5)>=5)), 5 , 0.01 ) }
 
 
** SWITCH 2 **
*
* ESD PROTECTION DIODES
D21 8 9 DCLAMP
D22 9 5 DCLAMP
D23 8 2 DCLAMP
D24 2 5 DCLAMP
*
* OFF ISOLATION
C21 2 9 1.9E-012
*
* CHARGE INJECTION
C22 9 240 2E-012
C23 2 240 2E-012
*
* CD/CS OFF AND BANDWIDTH
C24 2 4 12E-012
C25 9 4 15e-012
*
* ON RESISTANCE
Ech255 2555 4 VALUE = { IF ((ABS(V(2)))>(ABS(V(284))),V(2),V(9)) }
R255 2555 4 1G
R21 237 9 0.001
S221 236 241 2241 4 VON
Ech221 2241 4 VALUE = { IF (V(2555)<-13.5,5,0) }
Ech21 241 4 VALUE = { IF (V(2555)<-13.5,1.66666666666668E-02*(V(2555)--13.5)+2.45,0) }
S222 236 246 2246 4 VON
Ech222 2246 4 VALUE = { IF ((V(2555)>=-13.5) & (V(2555)<=13.5),5,0) }
Ech22 246 4 VALUE = { IF ((V(2555)>=-13.5) & (V(2555)<=13.5),((2.45-1.7)/((-13.5--0.796884641094606)*(-13.5--0.796884641094606)))*(V(2555)--0.796884641094606)*(V(2555)--0.796884641094606) + 1.7,0) }
S223 236 244 2244 4 VON
Ech223 2244 4 VALUE = { IF (V(2555)>13.5,5,0) }
Ech23 244 4 VALUE = { IF (V(2555)>13.5,-1.66666666666666E-02*(V(2555)-13.5)+2.65,0) }
RIN2	236 4	1G
EOUT2 237 281	POLY(2) (236,4) (280,4) 0 0 0 0 0.999/1000
FCOPY2	4 280 VSENSE2 1
RSENSOR2 280 4	1K
VSENSE2 281 284	0
*
* TON/ TOFF/ BBM
S21 282 284 240 4 VON
S22 243 238 243 4 VEN
Ech24 243 4 VALUE = { IF(V(6)>=2.0, 5 , 0.8 ) }
eV2 240 4 238 4 1
C26 238 4 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S23 2 282 285 4 VON
S24 242 285 242 4 VON
Ech25 242 4 VALUE = { IF((V(8)<=-0.5 & V(8)>=-16.5) & (V(5)<=16.5 & V(5)>=4.5), 5 , 0.01 ) }
S25 239 285 239 4 VON
Ech26 239 4 VALUE = { IF((V(8)>=-0.5 & (V(5)<=16.5 & V(5)>=5)), 5 , 0.01 ) }
 
.ENDS ADG1421
